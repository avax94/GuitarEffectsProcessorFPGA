library verilog;
use verilog.vl_types.all;
entity test_vibrato is
end test_vibrato;
