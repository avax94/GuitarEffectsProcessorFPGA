	// megafunction wizard: %SRAM/SSRAM Controller v13.0%
// GENERATION: XML
// sram.v

// Generated using ACDS version 13.0sp1 232 at 2018.05.01.15:33:39

`timescale 1 ps / 1 ps
module sram (
		input  wire        clk,           //        clock_reset.clk
		input  wire        reset,         //  clock_reset_reset.reset
		inout  wire [15:0] SRAM_DQ,       // external_interface.export
		output wire [17:0] SRAM_ADDR,     //                   .export
		output wire        SRAM_LB_N,     //                   .export
		output wire        SRAM_UB_N,     //                   .export
		output wire        SRAM_CE_N,     //                   .export
		output wire        SRAM_OE_N,     //                   .export
		output wire        SRAM_WE_N,     //                   .export
		input  wire [17:0] address,       //  avalon_sram_slave.address
		input  wire [1:0]  byteenable,    //                   .byteenable
		input  wire        read,          //                   .read
		input  wire        write,         //                   .write
		input  wire [15:0] writedata,     //                   .writedata
		output wire [15:0] readdata,      //                   .readdata
		output wire        readdatavalid  //                   .readdatavalid
	);

	sram_0002 sram_inst (
		.clk           (clk),           //        clock_reset.clk
		.reset         (reset),         //  clock_reset_reset.reset
		.SRAM_DQ       (SRAM_DQ),       // external_interface.export
		.SRAM_ADDR     (SRAM_ADDR),     //                   .export
		.SRAM_LB_N     (SRAM_LB_N),     //                   .export
		.SRAM_UB_N     (SRAM_UB_N),     //                   .export
		.SRAM_CE_N     (SRAM_CE_N),     //                   .export
		.SRAM_OE_N     (SRAM_OE_N),     //                   .export
		.SRAM_WE_N     (SRAM_WE_N),     //                   .export
		.address       (address),       //  avalon_sram_slave.address
		.byteenable    (byteenable),    //                   .byteenable
		.read          (read),          //                   .read
		.write         (write),         //                   .write
		.writedata     (writedata),     //                   .writedata
		.readdata      (readdata),      //                   .readdata
		.readdatavalid (readdatavalid)  //                   .readdatavalid
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2018 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_up_avalon_sram" version="13.0" >
// Retrieval info: 	<generic name="board" value="DE1" />
// Retrieval info: 	<generic name="pixel_buffer" value="false" />
// Retrieval info: 	<generic name="AUTO_CLOCK_RESET_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone II" />
// Retrieval info: </instance>
// IPFS_FILES : sram.vo
// RELATED_FILES: sram.v, sram_0002.v
