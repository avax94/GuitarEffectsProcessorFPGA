// megafunction wizard: %Audio and Video Config v13.0%
// GENERATION: XML
// av_config.v

// Generated using ACDS version 13.0sp1 232 at 2018.04.28.12:27:09

`timescale 1 ps / 1 ps
module av_config (
		input  wire        clk,         //            clock_reset.clk
		input  wire        reset,       //      clock_reset_reset.reset
		input  wire [1:0]  address,     // avalon_av_config_slave.address
		input  wire [3:0]  byteenable,  //                       .byteenable
		input  wire        read,        //                       .read
		input  wire        write,       //                       .write
		input  wire [31:0] writedata,   //                       .writedata
		output wire [31:0] readdata,    //                       .readdata
		output wire        waitrequest, //                       .waitrequest
		inout  wire        I2C_SDAT,    //     external_interface.export
		output wire        I2C_SCLK     //                       .export
	);

	av_config_0002 av_config_inst (
		.clk         (clk),         //            clock_reset.clk
		.reset       (reset),       //      clock_reset_reset.reset
		.address     (address),     // avalon_av_config_slave.address
		.byteenable  (byteenable),  //                       .byteenable
		.read        (read),        //                       .read
		.write       (write),       //                       .write
		.writedata   (writedata),   //                       .writedata
		.readdata    (readdata),    //                       .readdata
		.waitrequest (waitrequest), //                       .waitrequest
		.I2C_SDAT    (I2C_SDAT),    //     external_interface.export
		.I2C_SCLK    (I2C_SCLK)     //                       .export
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2018 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_up_avalon_audio_and_video_config" version="13.0" >
// Retrieval info: 	<generic name="device" value="On-Board Peripherals" />
// Retrieval info: 	<generic name="board" value="DE1" />
// Retrieval info: 	<generic name="eai" value="true" />
// Retrieval info: 	<generic name="audio_in" value="Microphone to ADC" />
// Retrieval info: 	<generic name="dac_enable" value="true" />
// Retrieval info: 	<generic name="mic_bypass" value="false" />
// Retrieval info: 	<generic name="line_in_bypass" value="false" />
// Retrieval info: 	<generic name="mic_attenuation" value="-6dB" />
// Retrieval info: 	<generic name="data_format" value="Left Justified" />
// Retrieval info: 	<generic name="bit_length" value="16" />
// Retrieval info: 	<generic name="sampling_rate" value="48 kHz" />
// Retrieval info: 	<generic name="video_format" value="NTSC" />
// Retrieval info: 	<generic name="d5m_resolution" value="2592 x 1944" />
// Retrieval info: 	<generic name="exposure" value="false" />
// Retrieval info: 	<generic name="AUTO_CLOCK_RESET_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone II" />
// Retrieval info: </instance>
// IPFS_FILES : av_config.vo
// RELATED_FILES: av_config.v, altera_up_av_config_serial_bus_controller.v, altera_up_slow_clock_generator.v, altera_up_av_config_auto_init.v, altera_up_av_config_auto_init_dc2.v, altera_up_av_config_auto_init_d5m.v, altera_up_av_config_auto_init_lcm.v, altera_up_av_config_auto_init_ltm.v, altera_up_av_config_auto_init_ob_de2_35.v, altera_up_av_config_auto_init_ob_adv7181.v, altera_up_av_config_auto_init_ob_de2_70.v, altera_up_av_config_auto_init_ob_de2_115.v, altera_up_av_config_auto_init_ob_audio.v, altera_up_av_config_auto_init_ob_adv7180.v, av_config_0002.v
