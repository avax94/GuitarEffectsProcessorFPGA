library verilog;
use verilog.vl_types.all;
entity test_smart_ram is
end test_smart_ram;
