library verilog;
use verilog.vl_types.all;
entity sinus_altfp_sincos_cordic_start_339 is
    port(
        index           : in     vl_logic_vector(3 downto 0);
        value           : out    vl_logic_vector(33 downto 0)
    );
end sinus_altfp_sincos_cordic_start_339;
