library verilog;
use verilog.vl_types.all;
entity test_noise_filter is
end test_noise_filter;
