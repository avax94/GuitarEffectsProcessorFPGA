// megafunction wizard: %Clock Signals for DE-series Board Peripherals v13.0%
// GENERATION: XML
// audio_clock_gen.v

// Generated using ACDS version 13.0sp1 232 at 2018.04.28.12:31:38

`timescale 1 ps / 1 ps
module audio_clock_gen (
		input  wire  CLOCK_50,    //       clk_in_primary.clk
		input  wire  reset,       // clk_in_primary_reset.reset
		output wire  sys_clk,     //              sys_clk.clk
		output wire  sys_reset_n, //        sys_clk_reset.reset_n
		output wire  SDRAM_CLK,   //            sdram_clk.clk
		input  wire  CLOCK_27,    //     clk_in_secondary.clk
		output wire  AUD_CLK      //            audio_clk.clk
	);

	audio_clock_gen_0002 audio_clock_gen_inst (
		.CLOCK_50    (CLOCK_50),    //       clk_in_primary.clk
		.reset       (reset),       // clk_in_primary_reset.reset
		.sys_clk     (sys_clk),     //              sys_clk.clk
		.sys_reset_n (sys_reset_n), //        sys_clk_reset.reset_n
		.SDRAM_CLK   (SDRAM_CLK),   //            sdram_clk.clk
		.CLOCK_27    (CLOCK_27),    //     clk_in_secondary.clk
		.AUD_CLK     (AUD_CLK)      //            audio_clk.clk
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2018 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_up_clocks" version="13.0" >
// Retrieval info: 	<generic name="board" value="DE1" />
// Retrieval info: 	<generic name="sys_clk_freq" value="50" />
// Retrieval info: 	<generic name="sdram_clk" value="true" />
// Retrieval info: 	<generic name="vga_clk" value="false" />
// Retrieval info: 	<generic name="audio_clk" value="true" />
// Retrieval info: 	<generic name="audio_clk_freq" value="12.288" />
// Retrieval info: 	<generic name="AUTO_CLK_IN_PRIMARY_CLOCK_RATE" value="-1" />
// Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone II" />
// Retrieval info: </instance>
// IPFS_FILES : audio_clock_gen.vo
// RELATED_FILES: audio_clock_gen.v, audio_clock_gen_0002.v
