library verilog;
use verilog.vl_types.all;
entity sinus_altpriority_encoder_0c6 is
    port(
        data            : in     vl_logic_vector(63 downto 0);
        q               : out    vl_logic_vector(5 downto 0)
    );
end sinus_altpriority_encoder_0c6;
