library verilog;
use verilog.vl_types.all;
entity test_echo is
end test_echo;
