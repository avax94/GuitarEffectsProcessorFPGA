library verilog;
use verilog.vl_types.all;
entity test_chorus is
end test_chorus;
